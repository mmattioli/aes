--
-- Written by Michael Mattioli
--
-- Description: AES package.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package aes is

    constant rounds : integer := 10; -- 10 rounds.

end aes;